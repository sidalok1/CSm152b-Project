`ifndef DEF_MAC
`define DEF_MAC

`define DATA_SIZE 8

`else

`endif
