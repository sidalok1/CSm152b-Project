$readmemh("k1_0-0.mem", conv1.kernels[0][0]);
$readmemh("k1_0-1.mem", conv1.kernels[0][1]);
$readmemh("k1_0-2.mem", conv1.kernels[0][2]);
$readmemh("k1_0-3.mem", conv1.kernels[0][3]);
$readmemh("k1_0-4.mem", conv1.kernels[0][4]);
$readmemh("k1_0-5.mem", conv1.kernels[0][5]);
$readmemh("k1_0-6.mem", conv1.kernels[0][6]);
$readmemh("k1_0-7.mem", conv1.kernels[0][7]);
$readmemh("k1_0-8.mem", conv1.kernels[0][8]);
$readmemh("k1_0-9.mem", conv1.kernels[0][9]);
$readmemh("k1_0-10.mem", conv1.kernels[0][10]);
$readmemh("k1_0-11.mem", conv1.kernels[0][11]);
$readmemh("k1_0-12.mem", conv1.kernels[0][12]);
$readmemh("k1_0-13.mem", conv1.kernels[0][13]);
$readmemh("k1_0-14.mem", conv1.kernels[0][14]);
$readmemh("k1_0-15.mem", conv1.kernels[0][15]);
$readmemh("k2_0-0.mem", conv2.kernels[0][0]);
$readmemh("k2_0-1.mem", conv2.kernels[0][1]);
$readmemh("k2_0-2.mem", conv2.kernels[0][2]);
$readmemh("k2_0-3.mem", conv2.kernels[0][3]);
$readmemh("k2_0-4.mem", conv2.kernels[0][4]);
$readmemh("k2_0-5.mem", conv2.kernels[0][5]);
$readmemh("k2_0-6.mem", conv2.kernels[0][6]);
$readmemh("k2_0-7.mem", conv2.kernels[0][7]);
$readmemh("k2_0-8.mem", conv2.kernels[0][8]);
$readmemh("k2_0-9.mem", conv2.kernels[0][9]);
$readmemh("k2_0-10.mem", conv2.kernels[0][10]);
$readmemh("k2_0-11.mem", conv2.kernels[0][11]);
$readmemh("k2_0-12.mem", conv2.kernels[0][12]);
$readmemh("k2_0-13.mem", conv2.kernels[0][13]);
$readmemh("k2_0-14.mem", conv2.kernels[0][14]);
$readmemh("k2_0-15.mem", conv2.kernels[0][15]);
$readmemh("k2_0-16.mem", conv2.kernels[0][16]);
$readmemh("k2_0-17.mem", conv2.kernels[0][17]);
$readmemh("k2_0-18.mem", conv2.kernels[0][18]);
$readmemh("k2_0-19.mem", conv2.kernels[0][19]);
$readmemh("k2_0-20.mem", conv2.kernels[0][20]);
$readmemh("k2_0-21.mem", conv2.kernels[0][21]);
$readmemh("k2_0-22.mem", conv2.kernels[0][22]);
$readmemh("k2_0-23.mem", conv2.kernels[0][23]);
$readmemh("k2_0-24.mem", conv2.kernels[0][24]);
$readmemh("k2_0-25.mem", conv2.kernels[0][25]);
$readmemh("k2_0-26.mem", conv2.kernels[0][26]);
$readmemh("k2_0-27.mem", conv2.kernels[0][27]);
$readmemh("k2_0-28.mem", conv2.kernels[0][28]);
$readmemh("k2_0-29.mem", conv2.kernels[0][29]);
$readmemh("k2_0-30.mem", conv2.kernels[0][30]);
$readmemh("k2_0-31.mem", conv2.kernels[0][31]);
$readmemh("k2_1-0.mem", conv2.kernels[1][0]);
$readmemh("k2_1-1.mem", conv2.kernels[1][1]);
$readmemh("k2_1-2.mem", conv2.kernels[1][2]);
$readmemh("k2_1-3.mem", conv2.kernels[1][3]);
$readmemh("k2_1-4.mem", conv2.kernels[1][4]);
$readmemh("k2_1-5.mem", conv2.kernels[1][5]);
$readmemh("k2_1-6.mem", conv2.kernels[1][6]);
$readmemh("k2_1-7.mem", conv2.kernels[1][7]);
$readmemh("k2_1-8.mem", conv2.kernels[1][8]);
$readmemh("k2_1-9.mem", conv2.kernels[1][9]);
$readmemh("k2_1-10.mem", conv2.kernels[1][10]);
$readmemh("k2_1-11.mem", conv2.kernels[1][11]);
$readmemh("k2_1-12.mem", conv2.kernels[1][12]);
$readmemh("k2_1-13.mem", conv2.kernels[1][13]);
$readmemh("k2_1-14.mem", conv2.kernels[1][14]);
$readmemh("k2_1-15.mem", conv2.kernels[1][15]);
$readmemh("k2_1-16.mem", conv2.kernels[1][16]);
$readmemh("k2_1-17.mem", conv2.kernels[1][17]);
$readmemh("k2_1-18.mem", conv2.kernels[1][18]);
$readmemh("k2_1-19.mem", conv2.kernels[1][19]);
$readmemh("k2_1-20.mem", conv2.kernels[1][20]);
$readmemh("k2_1-21.mem", conv2.kernels[1][21]);
$readmemh("k2_1-22.mem", conv2.kernels[1][22]);
$readmemh("k2_1-23.mem", conv2.kernels[1][23]);
$readmemh("k2_1-24.mem", conv2.kernels[1][24]);
$readmemh("k2_1-25.mem", conv2.kernels[1][25]);
$readmemh("k2_1-26.mem", conv2.kernels[1][26]);
$readmemh("k2_1-27.mem", conv2.kernels[1][27]);
$readmemh("k2_1-28.mem", conv2.kernels[1][28]);
$readmemh("k2_1-29.mem", conv2.kernels[1][29]);
$readmemh("k2_1-30.mem", conv2.kernels[1][30]);
$readmemh("k2_1-31.mem", conv2.kernels[1][31]);
$readmemh("k2_2-0.mem", conv2.kernels[2][0]);
$readmemh("k2_2-1.mem", conv2.kernels[2][1]);
$readmemh("k2_2-2.mem", conv2.kernels[2][2]);
$readmemh("k2_2-3.mem", conv2.kernels[2][3]);
$readmemh("k2_2-4.mem", conv2.kernels[2][4]);
$readmemh("k2_2-5.mem", conv2.kernels[2][5]);
$readmemh("k2_2-6.mem", conv2.kernels[2][6]);
$readmemh("k2_2-7.mem", conv2.kernels[2][7]);
$readmemh("k2_2-8.mem", conv2.kernels[2][8]);
$readmemh("k2_2-9.mem", conv2.kernels[2][9]);
$readmemh("k2_2-10.mem", conv2.kernels[2][10]);
$readmemh("k2_2-11.mem", conv2.kernels[2][11]);
$readmemh("k2_2-12.mem", conv2.kernels[2][12]);
$readmemh("k2_2-13.mem", conv2.kernels[2][13]);
$readmemh("k2_2-14.mem", conv2.kernels[2][14]);
$readmemh("k2_2-15.mem", conv2.kernels[2][15]);
$readmemh("k2_2-16.mem", conv2.kernels[2][16]);
$readmemh("k2_2-17.mem", conv2.kernels[2][17]);
$readmemh("k2_2-18.mem", conv2.kernels[2][18]);
$readmemh("k2_2-19.mem", conv2.kernels[2][19]);
$readmemh("k2_2-20.mem", conv2.kernels[2][20]);
$readmemh("k2_2-21.mem", conv2.kernels[2][21]);
$readmemh("k2_2-22.mem", conv2.kernels[2][22]);
$readmemh("k2_2-23.mem", conv2.kernels[2][23]);
$readmemh("k2_2-24.mem", conv2.kernels[2][24]);
$readmemh("k2_2-25.mem", conv2.kernels[2][25]);
$readmemh("k2_2-26.mem", conv2.kernels[2][26]);
$readmemh("k2_2-27.mem", conv2.kernels[2][27]);
$readmemh("k2_2-28.mem", conv2.kernels[2][28]);
$readmemh("k2_2-29.mem", conv2.kernels[2][29]);
$readmemh("k2_2-30.mem", conv2.kernels[2][30]);
$readmemh("k2_2-31.mem", conv2.kernels[2][31]);
$readmemh("k2_3-0.mem", conv2.kernels[3][0]);
$readmemh("k2_3-1.mem", conv2.kernels[3][1]);
$readmemh("k2_3-2.mem", conv2.kernels[3][2]);
$readmemh("k2_3-3.mem", conv2.kernels[3][3]);
$readmemh("k2_3-4.mem", conv2.kernels[3][4]);
$readmemh("k2_3-5.mem", conv2.kernels[3][5]);
$readmemh("k2_3-6.mem", conv2.kernels[3][6]);
$readmemh("k2_3-7.mem", conv2.kernels[3][7]);
$readmemh("k2_3-8.mem", conv2.kernels[3][8]);
$readmemh("k2_3-9.mem", conv2.kernels[3][9]);
$readmemh("k2_3-10.mem", conv2.kernels[3][10]);
$readmemh("k2_3-11.mem", conv2.kernels[3][11]);
$readmemh("k2_3-12.mem", conv2.kernels[3][12]);
$readmemh("k2_3-13.mem", conv2.kernels[3][13]);
$readmemh("k2_3-14.mem", conv2.kernels[3][14]);
$readmemh("k2_3-15.mem", conv2.kernels[3][15]);
$readmemh("k2_3-16.mem", conv2.kernels[3][16]);
$readmemh("k2_3-17.mem", conv2.kernels[3][17]);
$readmemh("k2_3-18.mem", conv2.kernels[3][18]);
$readmemh("k2_3-19.mem", conv2.kernels[3][19]);
$readmemh("k2_3-20.mem", conv2.kernels[3][20]);
$readmemh("k2_3-21.mem", conv2.kernels[3][21]);
$readmemh("k2_3-22.mem", conv2.kernels[3][22]);
$readmemh("k2_3-23.mem", conv2.kernels[3][23]);
$readmemh("k2_3-24.mem", conv2.kernels[3][24]);
$readmemh("k2_3-25.mem", conv2.kernels[3][25]);
$readmemh("k2_3-26.mem", conv2.kernels[3][26]);
$readmemh("k2_3-27.mem", conv2.kernels[3][27]);
$readmemh("k2_3-28.mem", conv2.kernels[3][28]);
$readmemh("k2_3-29.mem", conv2.kernels[3][29]);
$readmemh("k2_3-30.mem", conv2.kernels[3][30]);
$readmemh("k2_3-31.mem", conv2.kernels[3][31]);
$readmemh("k2_4-0.mem", conv2.kernels[4][0]);
$readmemh("k2_4-1.mem", conv2.kernels[4][1]);
$readmemh("k2_4-2.mem", conv2.kernels[4][2]);
$readmemh("k2_4-3.mem", conv2.kernels[4][3]);
$readmemh("k2_4-4.mem", conv2.kernels[4][4]);
$readmemh("k2_4-5.mem", conv2.kernels[4][5]);
$readmemh("k2_4-6.mem", conv2.kernels[4][6]);
$readmemh("k2_4-7.mem", conv2.kernels[4][7]);
$readmemh("k2_4-8.mem", conv2.kernels[4][8]);
$readmemh("k2_4-9.mem", conv2.kernels[4][9]);
$readmemh("k2_4-10.mem", conv2.kernels[4][10]);
$readmemh("k2_4-11.mem", conv2.kernels[4][11]);
$readmemh("k2_4-12.mem", conv2.kernels[4][12]);
$readmemh("k2_4-13.mem", conv2.kernels[4][13]);
$readmemh("k2_4-14.mem", conv2.kernels[4][14]);
$readmemh("k2_4-15.mem", conv2.kernels[4][15]);
$readmemh("k2_4-16.mem", conv2.kernels[4][16]);
$readmemh("k2_4-17.mem", conv2.kernels[4][17]);
$readmemh("k2_4-18.mem", conv2.kernels[4][18]);
$readmemh("k2_4-19.mem", conv2.kernels[4][19]);
$readmemh("k2_4-20.mem", conv2.kernels[4][20]);
$readmemh("k2_4-21.mem", conv2.kernels[4][21]);
$readmemh("k2_4-22.mem", conv2.kernels[4][22]);
$readmemh("k2_4-23.mem", conv2.kernels[4][23]);
$readmemh("k2_4-24.mem", conv2.kernels[4][24]);
$readmemh("k2_4-25.mem", conv2.kernels[4][25]);
$readmemh("k2_4-26.mem", conv2.kernels[4][26]);
$readmemh("k2_4-27.mem", conv2.kernels[4][27]);
$readmemh("k2_4-28.mem", conv2.kernels[4][28]);
$readmemh("k2_4-29.mem", conv2.kernels[4][29]);
$readmemh("k2_4-30.mem", conv2.kernels[4][30]);
$readmemh("k2_4-31.mem", conv2.kernels[4][31]);
$readmemh("k2_5-0.mem", conv2.kernels[5][0]);
$readmemh("k2_5-1.mem", conv2.kernels[5][1]);
$readmemh("k2_5-2.mem", conv2.kernels[5][2]);
$readmemh("k2_5-3.mem", conv2.kernels[5][3]);
$readmemh("k2_5-4.mem", conv2.kernels[5][4]);
$readmemh("k2_5-5.mem", conv2.kernels[5][5]);
$readmemh("k2_5-6.mem", conv2.kernels[5][6]);
$readmemh("k2_5-7.mem", conv2.kernels[5][7]);
$readmemh("k2_5-8.mem", conv2.kernels[5][8]);
$readmemh("k2_5-9.mem", conv2.kernels[5][9]);
$readmemh("k2_5-10.mem", conv2.kernels[5][10]);
$readmemh("k2_5-11.mem", conv2.kernels[5][11]);
$readmemh("k2_5-12.mem", conv2.kernels[5][12]);
$readmemh("k2_5-13.mem", conv2.kernels[5][13]);
$readmemh("k2_5-14.mem", conv2.kernels[5][14]);
$readmemh("k2_5-15.mem", conv2.kernels[5][15]);
$readmemh("k2_5-16.mem", conv2.kernels[5][16]);
$readmemh("k2_5-17.mem", conv2.kernels[5][17]);
$readmemh("k2_5-18.mem", conv2.kernels[5][18]);
$readmemh("k2_5-19.mem", conv2.kernels[5][19]);
$readmemh("k2_5-20.mem", conv2.kernels[5][20]);
$readmemh("k2_5-21.mem", conv2.kernels[5][21]);
$readmemh("k2_5-22.mem", conv2.kernels[5][22]);
$readmemh("k2_5-23.mem", conv2.kernels[5][23]);
$readmemh("k2_5-24.mem", conv2.kernels[5][24]);
$readmemh("k2_5-25.mem", conv2.kernels[5][25]);
$readmemh("k2_5-26.mem", conv2.kernels[5][26]);
$readmemh("k2_5-27.mem", conv2.kernels[5][27]);
$readmemh("k2_5-28.mem", conv2.kernels[5][28]);
$readmemh("k2_5-29.mem", conv2.kernels[5][29]);
$readmemh("k2_5-30.mem", conv2.kernels[5][30]);
$readmemh("k2_5-31.mem", conv2.kernels[5][31]);
$readmemh("k2_6-0.mem", conv2.kernels[6][0]);
$readmemh("k2_6-1.mem", conv2.kernels[6][1]);
$readmemh("k2_6-2.mem", conv2.kernels[6][2]);
$readmemh("k2_6-3.mem", conv2.kernels[6][3]);
$readmemh("k2_6-4.mem", conv2.kernels[6][4]);
$readmemh("k2_6-5.mem", conv2.kernels[6][5]);
$readmemh("k2_6-6.mem", conv2.kernels[6][6]);
$readmemh("k2_6-7.mem", conv2.kernels[6][7]);
$readmemh("k2_6-8.mem", conv2.kernels[6][8]);
$readmemh("k2_6-9.mem", conv2.kernels[6][9]);
$readmemh("k2_6-10.mem", conv2.kernels[6][10]);
$readmemh("k2_6-11.mem", conv2.kernels[6][11]);
$readmemh("k2_6-12.mem", conv2.kernels[6][12]);
$readmemh("k2_6-13.mem", conv2.kernels[6][13]);
$readmemh("k2_6-14.mem", conv2.kernels[6][14]);
$readmemh("k2_6-15.mem", conv2.kernels[6][15]);
$readmemh("k2_6-16.mem", conv2.kernels[6][16]);
$readmemh("k2_6-17.mem", conv2.kernels[6][17]);
$readmemh("k2_6-18.mem", conv2.kernels[6][18]);
$readmemh("k2_6-19.mem", conv2.kernels[6][19]);
$readmemh("k2_6-20.mem", conv2.kernels[6][20]);
$readmemh("k2_6-21.mem", conv2.kernels[6][21]);
$readmemh("k2_6-22.mem", conv2.kernels[6][22]);
$readmemh("k2_6-23.mem", conv2.kernels[6][23]);
$readmemh("k2_6-24.mem", conv2.kernels[6][24]);
$readmemh("k2_6-25.mem", conv2.kernels[6][25]);
$readmemh("k2_6-26.mem", conv2.kernels[6][26]);
$readmemh("k2_6-27.mem", conv2.kernels[6][27]);
$readmemh("k2_6-28.mem", conv2.kernels[6][28]);
$readmemh("k2_6-29.mem", conv2.kernels[6][29]);
$readmemh("k2_6-30.mem", conv2.kernels[6][30]);
$readmemh("k2_6-31.mem", conv2.kernels[6][31]);
$readmemh("k2_7-0.mem", conv2.kernels[7][0]);
$readmemh("k2_7-1.mem", conv2.kernels[7][1]);
$readmemh("k2_7-2.mem", conv2.kernels[7][2]);
$readmemh("k2_7-3.mem", conv2.kernels[7][3]);
$readmemh("k2_7-4.mem", conv2.kernels[7][4]);
$readmemh("k2_7-5.mem", conv2.kernels[7][5]);
$readmemh("k2_7-6.mem", conv2.kernels[7][6]);
$readmemh("k2_7-7.mem", conv2.kernels[7][7]);
$readmemh("k2_7-8.mem", conv2.kernels[7][8]);
$readmemh("k2_7-9.mem", conv2.kernels[7][9]);
$readmemh("k2_7-10.mem", conv2.kernels[7][10]);
$readmemh("k2_7-11.mem", conv2.kernels[7][11]);
$readmemh("k2_7-12.mem", conv2.kernels[7][12]);
$readmemh("k2_7-13.mem", conv2.kernels[7][13]);
$readmemh("k2_7-14.mem", conv2.kernels[7][14]);
$readmemh("k2_7-15.mem", conv2.kernels[7][15]);
$readmemh("k2_7-16.mem", conv2.kernels[7][16]);
$readmemh("k2_7-17.mem", conv2.kernels[7][17]);
$readmemh("k2_7-18.mem", conv2.kernels[7][18]);
$readmemh("k2_7-19.mem", conv2.kernels[7][19]);
$readmemh("k2_7-20.mem", conv2.kernels[7][20]);
$readmemh("k2_7-21.mem", conv2.kernels[7][21]);
$readmemh("k2_7-22.mem", conv2.kernels[7][22]);
$readmemh("k2_7-23.mem", conv2.kernels[7][23]);
$readmemh("k2_7-24.mem", conv2.kernels[7][24]);
$readmemh("k2_7-25.mem", conv2.kernels[7][25]);
$readmemh("k2_7-26.mem", conv2.kernels[7][26]);
$readmemh("k2_7-27.mem", conv2.kernels[7][27]);
$readmemh("k2_7-28.mem", conv2.kernels[7][28]);
$readmemh("k2_7-29.mem", conv2.kernels[7][29]);
$readmemh("k2_7-30.mem", conv2.kernels[7][30]);
$readmemh("k2_7-31.mem", conv2.kernels[7][31]);
$readmemh("k2_8-0.mem", conv2.kernels[8][0]);
$readmemh("k2_8-1.mem", conv2.kernels[8][1]);
$readmemh("k2_8-2.mem", conv2.kernels[8][2]);
$readmemh("k2_8-3.mem", conv2.kernels[8][3]);
$readmemh("k2_8-4.mem", conv2.kernels[8][4]);
$readmemh("k2_8-5.mem", conv2.kernels[8][5]);
$readmemh("k2_8-6.mem", conv2.kernels[8][6]);
$readmemh("k2_8-7.mem", conv2.kernels[8][7]);
$readmemh("k2_8-8.mem", conv2.kernels[8][8]);
$readmemh("k2_8-9.mem", conv2.kernels[8][9]);
$readmemh("k2_8-10.mem", conv2.kernels[8][10]);
$readmemh("k2_8-11.mem", conv2.kernels[8][11]);
$readmemh("k2_8-12.mem", conv2.kernels[8][12]);
$readmemh("k2_8-13.mem", conv2.kernels[8][13]);
$readmemh("k2_8-14.mem", conv2.kernels[8][14]);
$readmemh("k2_8-15.mem", conv2.kernels[8][15]);
$readmemh("k2_8-16.mem", conv2.kernels[8][16]);
$readmemh("k2_8-17.mem", conv2.kernels[8][17]);
$readmemh("k2_8-18.mem", conv2.kernels[8][18]);
$readmemh("k2_8-19.mem", conv2.kernels[8][19]);
$readmemh("k2_8-20.mem", conv2.kernels[8][20]);
$readmemh("k2_8-21.mem", conv2.kernels[8][21]);
$readmemh("k2_8-22.mem", conv2.kernels[8][22]);
$readmemh("k2_8-23.mem", conv2.kernels[8][23]);
$readmemh("k2_8-24.mem", conv2.kernels[8][24]);
$readmemh("k2_8-25.mem", conv2.kernels[8][25]);
$readmemh("k2_8-26.mem", conv2.kernels[8][26]);
$readmemh("k2_8-27.mem", conv2.kernels[8][27]);
$readmemh("k2_8-28.mem", conv2.kernels[8][28]);
$readmemh("k2_8-29.mem", conv2.kernels[8][29]);
$readmemh("k2_8-30.mem", conv2.kernels[8][30]);
$readmemh("k2_8-31.mem", conv2.kernels[8][31]);
$readmemh("k2_9-0.mem", conv2.kernels[9][0]);
$readmemh("k2_9-1.mem", conv2.kernels[9][1]);
$readmemh("k2_9-2.mem", conv2.kernels[9][2]);
$readmemh("k2_9-3.mem", conv2.kernels[9][3]);
$readmemh("k2_9-4.mem", conv2.kernels[9][4]);
$readmemh("k2_9-5.mem", conv2.kernels[9][5]);
$readmemh("k2_9-6.mem", conv2.kernels[9][6]);
$readmemh("k2_9-7.mem", conv2.kernels[9][7]);
$readmemh("k2_9-8.mem", conv2.kernels[9][8]);
$readmemh("k2_9-9.mem", conv2.kernels[9][9]);
$readmemh("k2_9-10.mem", conv2.kernels[9][10]);
$readmemh("k2_9-11.mem", conv2.kernels[9][11]);
$readmemh("k2_9-12.mem", conv2.kernels[9][12]);
$readmemh("k2_9-13.mem", conv2.kernels[9][13]);
$readmemh("k2_9-14.mem", conv2.kernels[9][14]);
$readmemh("k2_9-15.mem", conv2.kernels[9][15]);
$readmemh("k2_9-16.mem", conv2.kernels[9][16]);
$readmemh("k2_9-17.mem", conv2.kernels[9][17]);
$readmemh("k2_9-18.mem", conv2.kernels[9][18]);
$readmemh("k2_9-19.mem", conv2.kernels[9][19]);
$readmemh("k2_9-20.mem", conv2.kernels[9][20]);
$readmemh("k2_9-21.mem", conv2.kernels[9][21]);
$readmemh("k2_9-22.mem", conv2.kernels[9][22]);
$readmemh("k2_9-23.mem", conv2.kernels[9][23]);
$readmemh("k2_9-24.mem", conv2.kernels[9][24]);
$readmemh("k2_9-25.mem", conv2.kernels[9][25]);
$readmemh("k2_9-26.mem", conv2.kernels[9][26]);
$readmemh("k2_9-27.mem", conv2.kernels[9][27]);
$readmemh("k2_9-28.mem", conv2.kernels[9][28]);
$readmemh("k2_9-29.mem", conv2.kernels[9][29]);
$readmemh("k2_9-30.mem", conv2.kernels[9][30]);
$readmemh("k2_9-31.mem", conv2.kernels[9][31]);
$readmemh("k2_10-0.mem", conv2.kernels[10][0]);
$readmemh("k2_10-1.mem", conv2.kernels[10][1]);
$readmemh("k2_10-2.mem", conv2.kernels[10][2]);
$readmemh("k2_10-3.mem", conv2.kernels[10][3]);
$readmemh("k2_10-4.mem", conv2.kernels[10][4]);
$readmemh("k2_10-5.mem", conv2.kernels[10][5]);
$readmemh("k2_10-6.mem", conv2.kernels[10][6]);
$readmemh("k2_10-7.mem", conv2.kernels[10][7]);
$readmemh("k2_10-8.mem", conv2.kernels[10][8]);
$readmemh("k2_10-9.mem", conv2.kernels[10][9]);
$readmemh("k2_10-10.mem", conv2.kernels[10][10]);
$readmemh("k2_10-11.mem", conv2.kernels[10][11]);
$readmemh("k2_10-12.mem", conv2.kernels[10][12]);
$readmemh("k2_10-13.mem", conv2.kernels[10][13]);
$readmemh("k2_10-14.mem", conv2.kernels[10][14]);
$readmemh("k2_10-15.mem", conv2.kernels[10][15]);
$readmemh("k2_10-16.mem", conv2.kernels[10][16]);
$readmemh("k2_10-17.mem", conv2.kernels[10][17]);
$readmemh("k2_10-18.mem", conv2.kernels[10][18]);
$readmemh("k2_10-19.mem", conv2.kernels[10][19]);
$readmemh("k2_10-20.mem", conv2.kernels[10][20]);
$readmemh("k2_10-21.mem", conv2.kernels[10][21]);
$readmemh("k2_10-22.mem", conv2.kernels[10][22]);
$readmemh("k2_10-23.mem", conv2.kernels[10][23]);
$readmemh("k2_10-24.mem", conv2.kernels[10][24]);
$readmemh("k2_10-25.mem", conv2.kernels[10][25]);
$readmemh("k2_10-26.mem", conv2.kernels[10][26]);
$readmemh("k2_10-27.mem", conv2.kernels[10][27]);
$readmemh("k2_10-28.mem", conv2.kernels[10][28]);
$readmemh("k2_10-29.mem", conv2.kernels[10][29]);
$readmemh("k2_10-30.mem", conv2.kernels[10][30]);
$readmemh("k2_10-31.mem", conv2.kernels[10][31]);
$readmemh("k2_11-0.mem", conv2.kernels[11][0]);
$readmemh("k2_11-1.mem", conv2.kernels[11][1]);
$readmemh("k2_11-2.mem", conv2.kernels[11][2]);
$readmemh("k2_11-3.mem", conv2.kernels[11][3]);
$readmemh("k2_11-4.mem", conv2.kernels[11][4]);
$readmemh("k2_11-5.mem", conv2.kernels[11][5]);
$readmemh("k2_11-6.mem", conv2.kernels[11][6]);
$readmemh("k2_11-7.mem", conv2.kernels[11][7]);
$readmemh("k2_11-8.mem", conv2.kernels[11][8]);
$readmemh("k2_11-9.mem", conv2.kernels[11][9]);
$readmemh("k2_11-10.mem", conv2.kernels[11][10]);
$readmemh("k2_11-11.mem", conv2.kernels[11][11]);
$readmemh("k2_11-12.mem", conv2.kernels[11][12]);
$readmemh("k2_11-13.mem", conv2.kernels[11][13]);
$readmemh("k2_11-14.mem", conv2.kernels[11][14]);
$readmemh("k2_11-15.mem", conv2.kernels[11][15]);
$readmemh("k2_11-16.mem", conv2.kernels[11][16]);
$readmemh("k2_11-17.mem", conv2.kernels[11][17]);
$readmemh("k2_11-18.mem", conv2.kernels[11][18]);
$readmemh("k2_11-19.mem", conv2.kernels[11][19]);
$readmemh("k2_11-20.mem", conv2.kernels[11][20]);
$readmemh("k2_11-21.mem", conv2.kernels[11][21]);
$readmemh("k2_11-22.mem", conv2.kernels[11][22]);
$readmemh("k2_11-23.mem", conv2.kernels[11][23]);
$readmemh("k2_11-24.mem", conv2.kernels[11][24]);
$readmemh("k2_11-25.mem", conv2.kernels[11][25]);
$readmemh("k2_11-26.mem", conv2.kernels[11][26]);
$readmemh("k2_11-27.mem", conv2.kernels[11][27]);
$readmemh("k2_11-28.mem", conv2.kernels[11][28]);
$readmemh("k2_11-29.mem", conv2.kernels[11][29]);
$readmemh("k2_11-30.mem", conv2.kernels[11][30]);
$readmemh("k2_11-31.mem", conv2.kernels[11][31]);
$readmemh("k2_12-0.mem", conv2.kernels[12][0]);
$readmemh("k2_12-1.mem", conv2.kernels[12][1]);
$readmemh("k2_12-2.mem", conv2.kernels[12][2]);
$readmemh("k2_12-3.mem", conv2.kernels[12][3]);
$readmemh("k2_12-4.mem", conv2.kernels[12][4]);
$readmemh("k2_12-5.mem", conv2.kernels[12][5]);
$readmemh("k2_12-6.mem", conv2.kernels[12][6]);
$readmemh("k2_12-7.mem", conv2.kernels[12][7]);
$readmemh("k2_12-8.mem", conv2.kernels[12][8]);
$readmemh("k2_12-9.mem", conv2.kernels[12][9]);
$readmemh("k2_12-10.mem", conv2.kernels[12][10]);
$readmemh("k2_12-11.mem", conv2.kernels[12][11]);
$readmemh("k2_12-12.mem", conv2.kernels[12][12]);
$readmemh("k2_12-13.mem", conv2.kernels[12][13]);
$readmemh("k2_12-14.mem", conv2.kernels[12][14]);
$readmemh("k2_12-15.mem", conv2.kernels[12][15]);
$readmemh("k2_12-16.mem", conv2.kernels[12][16]);
$readmemh("k2_12-17.mem", conv2.kernels[12][17]);
$readmemh("k2_12-18.mem", conv2.kernels[12][18]);
$readmemh("k2_12-19.mem", conv2.kernels[12][19]);
$readmemh("k2_12-20.mem", conv2.kernels[12][20]);
$readmemh("k2_12-21.mem", conv2.kernels[12][21]);
$readmemh("k2_12-22.mem", conv2.kernels[12][22]);
$readmemh("k2_12-23.mem", conv2.kernels[12][23]);
$readmemh("k2_12-24.mem", conv2.kernels[12][24]);
$readmemh("k2_12-25.mem", conv2.kernels[12][25]);
$readmemh("k2_12-26.mem", conv2.kernels[12][26]);
$readmemh("k2_12-27.mem", conv2.kernels[12][27]);
$readmemh("k2_12-28.mem", conv2.kernels[12][28]);
$readmemh("k2_12-29.mem", conv2.kernels[12][29]);
$readmemh("k2_12-30.mem", conv2.kernels[12][30]);
$readmemh("k2_12-31.mem", conv2.kernels[12][31]);
$readmemh("k2_13-0.mem", conv2.kernels[13][0]);
$readmemh("k2_13-1.mem", conv2.kernels[13][1]);
$readmemh("k2_13-2.mem", conv2.kernels[13][2]);
$readmemh("k2_13-3.mem", conv2.kernels[13][3]);
$readmemh("k2_13-4.mem", conv2.kernels[13][4]);
$readmemh("k2_13-5.mem", conv2.kernels[13][5]);
$readmemh("k2_13-6.mem", conv2.kernels[13][6]);
$readmemh("k2_13-7.mem", conv2.kernels[13][7]);
$readmemh("k2_13-8.mem", conv2.kernels[13][8]);
$readmemh("k2_13-9.mem", conv2.kernels[13][9]);
$readmemh("k2_13-10.mem", conv2.kernels[13][10]);
$readmemh("k2_13-11.mem", conv2.kernels[13][11]);
$readmemh("k2_13-12.mem", conv2.kernels[13][12]);
$readmemh("k2_13-13.mem", conv2.kernels[13][13]);
$readmemh("k2_13-14.mem", conv2.kernels[13][14]);
$readmemh("k2_13-15.mem", conv2.kernels[13][15]);
$readmemh("k2_13-16.mem", conv2.kernels[13][16]);
$readmemh("k2_13-17.mem", conv2.kernels[13][17]);
$readmemh("k2_13-18.mem", conv2.kernels[13][18]);
$readmemh("k2_13-19.mem", conv2.kernels[13][19]);
$readmemh("k2_13-20.mem", conv2.kernels[13][20]);
$readmemh("k2_13-21.mem", conv2.kernels[13][21]);
$readmemh("k2_13-22.mem", conv2.kernels[13][22]);
$readmemh("k2_13-23.mem", conv2.kernels[13][23]);
$readmemh("k2_13-24.mem", conv2.kernels[13][24]);
$readmemh("k2_13-25.mem", conv2.kernels[13][25]);
$readmemh("k2_13-26.mem", conv2.kernels[13][26]);
$readmemh("k2_13-27.mem", conv2.kernels[13][27]);
$readmemh("k2_13-28.mem", conv2.kernels[13][28]);
$readmemh("k2_13-29.mem", conv2.kernels[13][29]);
$readmemh("k2_13-30.mem", conv2.kernels[13][30]);
$readmemh("k2_13-31.mem", conv2.kernels[13][31]);
$readmemh("k2_14-0.mem", conv2.kernels[14][0]);
$readmemh("k2_14-1.mem", conv2.kernels[14][1]);
$readmemh("k2_14-2.mem", conv2.kernels[14][2]);
$readmemh("k2_14-3.mem", conv2.kernels[14][3]);
$readmemh("k2_14-4.mem", conv2.kernels[14][4]);
$readmemh("k2_14-5.mem", conv2.kernels[14][5]);
$readmemh("k2_14-6.mem", conv2.kernels[14][6]);
$readmemh("k2_14-7.mem", conv2.kernels[14][7]);
$readmemh("k2_14-8.mem", conv2.kernels[14][8]);
$readmemh("k2_14-9.mem", conv2.kernels[14][9]);
$readmemh("k2_14-10.mem", conv2.kernels[14][10]);
$readmemh("k2_14-11.mem", conv2.kernels[14][11]);
$readmemh("k2_14-12.mem", conv2.kernels[14][12]);
$readmemh("k2_14-13.mem", conv2.kernels[14][13]);
$readmemh("k2_14-14.mem", conv2.kernels[14][14]);
$readmemh("k2_14-15.mem", conv2.kernels[14][15]);
$readmemh("k2_14-16.mem", conv2.kernels[14][16]);
$readmemh("k2_14-17.mem", conv2.kernels[14][17]);
$readmemh("k2_14-18.mem", conv2.kernels[14][18]);
$readmemh("k2_14-19.mem", conv2.kernels[14][19]);
$readmemh("k2_14-20.mem", conv2.kernels[14][20]);
$readmemh("k2_14-21.mem", conv2.kernels[14][21]);
$readmemh("k2_14-22.mem", conv2.kernels[14][22]);
$readmemh("k2_14-23.mem", conv2.kernels[14][23]);
$readmemh("k2_14-24.mem", conv2.kernels[14][24]);
$readmemh("k2_14-25.mem", conv2.kernels[14][25]);
$readmemh("k2_14-26.mem", conv2.kernels[14][26]);
$readmemh("k2_14-27.mem", conv2.kernels[14][27]);
$readmemh("k2_14-28.mem", conv2.kernels[14][28]);
$readmemh("k2_14-29.mem", conv2.kernels[14][29]);
$readmemh("k2_14-30.mem", conv2.kernels[14][30]);
$readmemh("k2_14-31.mem", conv2.kernels[14][31]);
$readmemh("k2_15-0.mem", conv2.kernels[15][0]);
$readmemh("k2_15-1.mem", conv2.kernels[15][1]);
$readmemh("k2_15-2.mem", conv2.kernels[15][2]);
$readmemh("k2_15-3.mem", conv2.kernels[15][3]);
$readmemh("k2_15-4.mem", conv2.kernels[15][4]);
$readmemh("k2_15-5.mem", conv2.kernels[15][5]);
$readmemh("k2_15-6.mem", conv2.kernels[15][6]);
$readmemh("k2_15-7.mem", conv2.kernels[15][7]);
$readmemh("k2_15-8.mem", conv2.kernels[15][8]);
$readmemh("k2_15-9.mem", conv2.kernels[15][9]);
$readmemh("k2_15-10.mem", conv2.kernels[15][10]);
$readmemh("k2_15-11.mem", conv2.kernels[15][11]);
$readmemh("k2_15-12.mem", conv2.kernels[15][12]);
$readmemh("k2_15-13.mem", conv2.kernels[15][13]);
$readmemh("k2_15-14.mem", conv2.kernels[15][14]);
$readmemh("k2_15-15.mem", conv2.kernels[15][15]);
$readmemh("k2_15-16.mem", conv2.kernels[15][16]);
$readmemh("k2_15-17.mem", conv2.kernels[15][17]);
$readmemh("k2_15-18.mem", conv2.kernels[15][18]);
$readmemh("k2_15-19.mem", conv2.kernels[15][19]);
$readmemh("k2_15-20.mem", conv2.kernels[15][20]);
$readmemh("k2_15-21.mem", conv2.kernels[15][21]);
$readmemh("k2_15-22.mem", conv2.kernels[15][22]);
$readmemh("k2_15-23.mem", conv2.kernels[15][23]);
$readmemh("k2_15-24.mem", conv2.kernels[15][24]);
$readmemh("k2_15-25.mem", conv2.kernels[15][25]);
$readmemh("k2_15-26.mem", conv2.kernels[15][26]);
$readmemh("k2_15-27.mem", conv2.kernels[15][27]);
$readmemh("k2_15-28.mem", conv2.kernels[15][28]);
$readmemh("k2_15-29.mem", conv2.kernels[15][29]);
$readmemh("k2_15-30.mem", conv2.kernels[15][30]);
$readmemh("k2_15-31.mem", conv2.kernels[15][31]);